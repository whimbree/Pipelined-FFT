library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package user_pkg is

constant DATA_WIDTH : positive := 32;
subtype DATA_RANGE is natural range DATA_WIDTH - 1 downto 0;

constant NUM_POINTS : positive := 1024;

type TWIDDLE_ARRAY is array (natural range <>) of std_logic_vector(DATA_RANGE);
subtype TWIDDLE_RANGE is natural range 0 to NUM_POINTS - 1;

constant TWIDDLE_FACTORS_REAL : TWIDDLE_ARRAY(TWIDDLE_RANGE) := (0 => x"7fffffff",1 => x"7fff6215",2 => x"7ffd8859",3 => x"7ffa72d1",4 => x"7ff62182",5 => x"7ff09477",6 => x"7fe9cbbf",7 => x"7fe1c76b",8 => x"7fd8878d",9 => x"7fce0c3e",
10 => x"7fc25596",11 => x"7fb563b2",12 => x"7fa736b4",13 => x"7f97cebc",14 => x"7f872bf2",15 => x"7f754e7f",16 => x"7f62368f",17 => x"7f4de450",18 => x"7f3857f5",19 => x"7f2191b3",
20 => x"7f0991c3",21 => x"7ef0585f",22 => x"7ed5e5c6",23 => x"7eba3a39",24 => x"7e9d55fc",25 => x"7e7f3956",26 => x"7e5fe493",27 => x"7e3f57fe",28 => x"7e1d93e9",29 => x"7dfa98a7",
30 => x"7dd6668e",31 => x"7db0fdf7",32 => x"7d8a5f3f",33 => x"7d628ac5",34 => x"7d3980ec",35 => x"7d0f4217",36 => x"7ce3ceb1",37 => x"7cb72724",38 => x"7c894bdd",39 => x"7c5a3d4f",
40 => x"7c29fbee",41 => x"7bf88830",42 => x"7bc5e28f",43 => x"7b920b89",44 => x"7b5d039d",45 => x"7b26cb4f",46 => x"7aef6323",47 => x"7ab6cba3",48 => x"7a7d055b",49 => x"7a4210d8",
50 => x"7a05eead",51 => x"79c89f6d",52 => x"798a23b1",53 => x"794a7c11",54 => x"7909a92c",55 => x"78c7aba1",56 => x"78848413",57 => x"78403328",58 => x"77fab988",59 => x"77b417df",
60 => x"776c4edb",61 => x"77235f2d",62 => x"76d94988",63 => x"768e0ea5",64 => x"7641af3c",65 => x"75f42c0a",66 => x"75a585cf",67 => x"7555bd4b",68 => x"7504d345",69 => x"74b2c883",
70 => x"745f9dd0",71 => x"740b53fa",72 => x"73b5ebd0",73 => x"735f6626",74 => x"7307c3cf",75 => x"72af05a6",76 => x"72552c84",77 => x"71fa3948",78 => x"719e2cd2",79 => x"71410804",
80 => x"70e2cbc6",81 => x"708378fe",82 => x"70231099",83 => x"6fc19385",84 => x"6f5f02b1",85 => x"6efb5f12",86 => x"6e96a99c",87 => x"6e30e349",88 => x"6dca0d14",89 => x"6d6227fa",
90 => x"6cf934fb",91 => x"6c8f351c",92 => x"6c242960",93 => x"6bb812d0",94 => x"6b4af278",95 => x"6adcc964",96 => x"6a6d98a4",97 => x"69fd614a",98 => x"698c246c",99 => x"6919e320",
100 => x"68a69e81",101 => x"683257aa",102 => x"67bd0fbc",103 => x"6746c7d7",104 => x"66cf811f",105 => x"66573cbb",106 => x"65ddfbd3",107 => x"6563bf92",108 => x"64e88926",109 => x"646c59bf",
110 => x"63ef328f",111 => x"637114cc",112 => x"62f201ac",113 => x"6271fa69",114 => x"61f1003e",115 => x"616f146b",116 => x"60ec382f",117 => x"60686cce",118 => x"5fe3b38d",119 => x"5f5e0db3",
120 => x"5ed77c89",121 => x"5e50015d",122 => x"5dc79d7c",123 => x"5d3e5236",124 => x"5cb420df",125 => x"5c290acc",126 => x"5b9d1153",127 => x"5b1035cf",128 => x"5a827999",129 => x"59f3de12",
130 => x"59646497",131 => x"58d40e8c",132 => x"5842dd54",133 => x"57b0d256",134 => x"571deef9",135 => x"568a34a9",136 => x"55f5a4d2",137 => x"556040e2",138 => x"54ca0a4a",139 => x"5433027d",
140 => x"539b2aef",141 => x"53028517",142 => x"5269126e",143 => x"51ced46e",144 => x"5133cc94",145 => x"5097fc5e",146 => x"4ffb654d",147 => x"4f5e08e3",148 => x"4ebfe8a4",149 => x"4e210617",
150 => x"4d8162c4",151 => x"4ce10034",152 => x"4c3fdff3",153 => x"4b9e038f",154 => x"4afb6c97",155 => x"4a581c9d",156 => x"49b41533",157 => x"490f57ee",158 => x"4869e664",159 => x"47c3c22e",
160 => x"471cece6",161 => x"46756827",162 => x"45cd358f",163 => x"452456bc",164 => x"447acd50",165 => x"43d09aec",166 => x"4325c135",167 => x"427a41d0",168 => x"41ce1e64",169 => x"4121589a",
170 => x"4073f21d",171 => x"3fc5ec97",172 => x"3f1749b7",173 => x"3e680b2c",174 => x"3db832a5",175 => x"3d07c1d5",176 => x"3c56ba70",177 => x"3ba51e29",178 => x"3af2eeb7",179 => x"3a402dd1",
180 => x"398cdd32",181 => x"38d8fe93",182 => x"382493b0",183 => x"376f9e46",184 => x"36ba2013",185 => x"36041ad8",186 => x"354d9056",187 => x"3496824f",188 => x"33def287",189 => x"3326e2c2",
190 => x"326e54c7",191 => x"31b54a5d",192 => x"30fbc54d",193 => x"3041c760",194 => x"2f875262",195 => x"2ecc681e",196 => x"2e110a61",197 => x"2d553afb",198 => x"2c98fbba",199 => x"2bdc4e6f",
200 => x"2b1f34eb",201 => x"2a61b101",202 => x"29a3c484",203 => x"28e5714a",204 => x"2826b928",205 => x"27679df4",206 => x"26a82185",207 => x"25e845b5",208 => x"25280c5d",209 => x"24677757",
210 => x"23a6887e",211 => x"22e541ae",212 => x"2223a4c5",213 => x"2161b39f",214 => x"209f701c",215 => x"1fdcdc1a",216 => x"1f19f97b",217 => x"1e56ca1e",218 => x"1d934fe5",219 => x"1ccf8cb3",
220 => x"1c0b826a",221 => x"1b4732ef",222 => x"1a82a025",223 => x"19bdcbf2",224 => x"18f8b83c",225 => x"183366e8",226 => x"176dd9de",227 => x"16a81304",228 => x"15e21444",229 => x"151bdf85",
230 => x"145576b1",231 => x"138edbb0",232 => x"12c8106e",233 => x"120116d4",234 => x"1139f0ce",235 => x"1072a047",236 => x"0fab272b",237 => x"0ee38765",238 => x"0e1bc2e3",239 => x"0d53db92",
240 => x"0c8bd35e",241 => x"0bc3ac35",242 => x"0afb6805",243 => x"0a3308bc",244 => x"096a9049",245 => x"08a2009a",246 => x"07d95b9e",247 => x"0710a344",248 => x"0647d97c",249 => x"057f0034",
250 => x"04b6195d",251 => x"03ed26e6",252 => x"03242abe",253 => x"025b26d7",254 => x"01921d1f",255 => x"00c90f87",256 => x"00000000",257 => x"ff36f079",258 => x"fe6de2e1",259 => x"fda4d929",
260 => x"fcdbd542",261 => x"fc12d91a",262 => x"fb49e6a3",263 => x"fa80ffcc",264 => x"f9b82684",265 => x"f8ef5cbc",266 => x"f826a462",267 => x"f75dff66",268 => x"f6956fb7",269 => x"f5ccf744",
270 => x"f50497fb",271 => x"f43c53cb",272 => x"f3742ca2",273 => x"f2ac246e",274 => x"f1e43d1d",275 => x"f11c789b",276 => x"f054d8d5",277 => x"ef8d5fb9",278 => x"eec60f32",279 => x"edfee92c",
280 => x"ed37ef92",281 => x"ec712450",282 => x"ebaa894f",283 => x"eae4207b",284 => x"ea1debbc",285 => x"e957ecfc",286 => x"e8922622",287 => x"e7cc9918",288 => x"e70747c4",289 => x"e642340e",
290 => x"e57d5fdb",291 => x"e4b8cd11",292 => x"e3f47d96",293 => x"e330734d",294 => x"e26cb01b",295 => x"e1a935e2",296 => x"e0e60685",297 => x"e02323e6",298 => x"df608fe4",299 => x"de9e4c61",
300 => x"dddc5b3b",301 => x"dd1abe52",302 => x"dc597782",303 => x"db9888a9",304 => x"dad7f3a3",305 => x"da17ba4b",306 => x"d957de7b",307 => x"d898620c",308 => x"d7d946d8",309 => x"d71a8eb6",
310 => x"d65c3b7c",311 => x"d59e4eff",312 => x"d4e0cb15",313 => x"d423b191",314 => x"d3670446",315 => x"d2aac505",316 => x"d1eef59f",317 => x"d13397e2",318 => x"d078ad9e",319 => x"cfbe38a0",
320 => x"cf043ab3",321 => x"ce4ab5a3",322 => x"cd91ab39",323 => x"ccd91d3e",324 => x"cc210d79",325 => x"cb697db1",326 => x"cab26faa",327 => x"c9fbe528",328 => x"c945dfed",329 => x"c89061ba",
330 => x"c7db6c50",331 => x"c727016d",332 => x"c67322ce",333 => x"c5bfd22f",334 => x"c50d1149",335 => x"c45ae1d7",336 => x"c3a94590",337 => x"c2f83e2b",338 => x"c247cd5b",339 => x"c197f4d4",
340 => x"c0e8b649",341 => x"c03a1369",342 => x"bf8c0de3",343 => x"bedea766",344 => x"be31e19c",345 => x"bd85be30",346 => x"bcda3ecb",347 => x"bc2f6514",348 => x"bb8532b0",349 => x"badba944",
350 => x"ba32ca71",351 => x"b98a97d9",352 => x"b8e3131a",353 => x"b83c3dd2",354 => x"b796199c",355 => x"b6f0a812",356 => x"b64beacd",357 => x"b5a7e363",358 => x"b5049369",359 => x"b461fc71",
360 => x"b3c0200d",361 => x"b31effcc",362 => x"b27e9d3c",363 => x"b1def9e9",364 => x"b140175c",365 => x"b0a1f71d",366 => x"b0049ab3",367 => x"af6803a2",368 => x"aecc336c",369 => x"ae312b92",
370 => x"ad96ed92",371 => x"acfd7ae9",372 => x"ac64d511",373 => x"abccfd83",374 => x"ab35f5b6",375 => x"aa9fbf1e",376 => x"aa0a5b2e",377 => x"a975cb57",378 => x"a8e21107",379 => x"a84f2daa",
380 => x"a7bd22ac",381 => x"a72bf174",382 => x"a69b9b69",383 => x"a60c21ee",384 => x"a57d8667",385 => x"a4efca31",386 => x"a462eead",387 => x"a3d6f534",388 => x"a34bdf21",389 => x"a2c1adca",
390 => x"a2386284",391 => x"a1affea3",392 => x"a1288377",393 => x"a0a1f24d",394 => x"a01c4c73",395 => x"9f979332",396 => x"9f13c7d1",397 => x"9e90eb95",398 => x"9e0effc2",399 => x"9d8e0597",
400 => x"9d0dfe54",401 => x"9c8eeb34",402 => x"9c10cd71",403 => x"9b93a641",404 => x"9b1776da",405 => x"9a9c406e",406 => x"9a22042d",407 => x"99a8c345",408 => x"99307ee1",409 => x"98b93829",
410 => x"9842f044",411 => x"97cda856",412 => x"9759617f",413 => x"96e61ce0",414 => x"9673db94",415 => x"96029eb6",416 => x"9592675c",417 => x"9523369c",418 => x"94b50d88",419 => x"9447ed30",
420 => x"93dbd6a0",421 => x"9370cae4",422 => x"9306cb05",423 => x"929dd806",424 => x"9235f2ec",425 => x"91cf1cb7",426 => x"91695664",427 => x"9104a0ee",428 => x"90a0fd4f",429 => x"903e6c7b",
430 => x"8fdcef67",431 => x"8f7c8702",432 => x"8f1d343a",433 => x"8ebef7fc",434 => x"8e61d32e",435 => x"8e05c6b8",436 => x"8daad37c",437 => x"8d50fa5a",438 => x"8cf83c31",439 => x"8ca099da",
440 => x"8c4a1430",441 => x"8bf4ac06",442 => x"8ba06230",443 => x"8b4d377d",444 => x"8afb2cbb",445 => x"8aaa42b5",446 => x"8a5a7a31",447 => x"8a0bd3f6",448 => x"89be50c4",449 => x"8971f15b",
450 => x"8926b678",451 => x"88dca0d3",452 => x"8893b125",453 => x"884be821",454 => x"88054678",455 => x"87bfccd8",456 => x"877b7bed",457 => x"8738545f",458 => x"86f656d4",459 => x"86b583ef",
460 => x"8675dc4f",461 => x"86376093",462 => x"85fa1153",463 => x"85bdef28",464 => x"8582faa5",465 => x"8549345d",466 => x"85109cdd",467 => x"84d934b1",468 => x"84a2fc63",469 => x"846df477",
470 => x"843a1d71",471 => x"840777d0",472 => x"83d60412",473 => x"83a5c2b1",474 => x"8376b423",475 => x"8348d8dc",476 => x"831c314f",477 => x"82f0bde9",478 => x"82c67f14",479 => x"829d753b",
480 => x"8275a0c1",481 => x"824f0209",482 => x"82299972",483 => x"82056759",484 => x"81e26c17",485 => x"81c0a802",486 => x"81a01b6d",487 => x"8180c6aa",488 => x"8162aa04",489 => x"8145c5c7",
490 => x"812a1a3a",491 => x"810fa7a1",492 => x"80f66e3d",493 => x"80de6e4d",494 => x"80c7a80b",495 => x"80b21bb0",496 => x"809dc971",497 => x"808ab181",498 => x"8078d40e",499 => x"80683144",
500 => x"8058c94c",501 => x"804a9c4e",502 => x"803daa6a",503 => x"8031f3c2",504 => x"80277873",505 => x"801e3895",506 => x"80163441",507 => x"800f6b89",508 => x"8009de7e",509 => x"80058d2f",
510 => x"800277a6",511 => x"80009dea",512 => x"80000000",513 => x"80009dea",514 => x"800277a6",515 => x"80058d2f",516 => x"8009de7e",517 => x"800f6b89",518 => x"80163441",519 => x"801e3895",
520 => x"80277873",521 => x"8031f3c2",522 => x"803daa6a",523 => x"804a9c4e",524 => x"8058c94c",525 => x"80683144",526 => x"8078d40e",527 => x"808ab181",528 => x"809dc971",529 => x"80b21bb0",
530 => x"80c7a80b",531 => x"80de6e4d",532 => x"80f66e3d",533 => x"810fa7a1",534 => x"812a1a3a",535 => x"8145c5c7",536 => x"8162aa04",537 => x"8180c6aa",538 => x"81a01b6d",539 => x"81c0a802",
540 => x"81e26c17",541 => x"82056759",542 => x"82299972",543 => x"824f0209",544 => x"8275a0c1",545 => x"829d753b",546 => x"82c67f14",547 => x"82f0bde9",548 => x"831c314f",549 => x"8348d8dc",
550 => x"8376b423",551 => x"83a5c2b1",552 => x"83d60412",553 => x"840777d0",554 => x"843a1d71",555 => x"846df477",556 => x"84a2fc63",557 => x"84d934b1",558 => x"85109cdd",559 => x"8549345d",
560 => x"8582faa5",561 => x"85bdef28",562 => x"85fa1153",563 => x"86376093",564 => x"8675dc4f",565 => x"86b583ef",566 => x"86f656d4",567 => x"8738545f",568 => x"877b7bed",569 => x"87bfccd8",
570 => x"88054678",571 => x"884be821",572 => x"8893b125",573 => x"88dca0d3",574 => x"8926b678",575 => x"8971f15b",576 => x"89be50c4",577 => x"8a0bd3f6",578 => x"8a5a7a31",579 => x"8aaa42b5",
580 => x"8afb2cbb",581 => x"8b4d377d",582 => x"8ba06230",583 => x"8bf4ac06",584 => x"8c4a1430",585 => x"8ca099da",586 => x"8cf83c31",587 => x"8d50fa5a",588 => x"8daad37c",589 => x"8e05c6b8",
590 => x"8e61d32e",591 => x"8ebef7fc",592 => x"8f1d343a",593 => x"8f7c8702",594 => x"8fdcef67",595 => x"903e6c7b",596 => x"90a0fd4f",597 => x"9104a0ee",598 => x"91695664",599 => x"91cf1cb7",
600 => x"9235f2ec",601 => x"929dd806",602 => x"9306cb05",603 => x"9370cae4",604 => x"93dbd6a0",605 => x"9447ed30",606 => x"94b50d88",607 => x"9523369c",608 => x"9592675c",609 => x"96029eb6",
610 => x"9673db94",611 => x"96e61ce0",612 => x"9759617f",613 => x"97cda856",614 => x"9842f044",615 => x"98b93829",616 => x"99307ee1",617 => x"99a8c345",618 => x"9a22042d",619 => x"9a9c406e",
620 => x"9b1776da",621 => x"9b93a641",622 => x"9c10cd71",623 => x"9c8eeb34",624 => x"9d0dfe54",625 => x"9d8e0597",626 => x"9e0effc2",627 => x"9e90eb95",628 => x"9f13c7d1",629 => x"9f979332",
630 => x"a01c4c73",631 => x"a0a1f24d",632 => x"a1288377",633 => x"a1affea3",634 => x"a2386284",635 => x"a2c1adca",636 => x"a34bdf21",637 => x"a3d6f534",638 => x"a462eead",639 => x"a4efca31",
640 => x"a57d8667",641 => x"a60c21ee",642 => x"a69b9b69",643 => x"a72bf174",644 => x"a7bd22ac",645 => x"a84f2daa",646 => x"a8e21107",647 => x"a975cb57",648 => x"aa0a5b2e",649 => x"aa9fbf1e",
650 => x"ab35f5b6",651 => x"abccfd83",652 => x"ac64d511",653 => x"acfd7ae9",654 => x"ad96ed92",655 => x"ae312b92",656 => x"aecc336c",657 => x"af6803a2",658 => x"b0049ab3",659 => x"b0a1f71d",
660 => x"b140175c",661 => x"b1def9e9",662 => x"b27e9d3c",663 => x"b31effcc",664 => x"b3c0200d",665 => x"b461fc71",666 => x"b5049369",667 => x"b5a7e363",668 => x"b64beacd",669 => x"b6f0a812",
670 => x"b796199c",671 => x"b83c3dd2",672 => x"b8e3131a",673 => x"b98a97d9",674 => x"ba32ca71",675 => x"badba944",676 => x"bb8532b0",677 => x"bc2f6514",678 => x"bcda3ecb",679 => x"bd85be30",
680 => x"be31e19c",681 => x"bedea766",682 => x"bf8c0de3",683 => x"c03a1369",684 => x"c0e8b649",685 => x"c197f4d4",686 => x"c247cd5b",687 => x"c2f83e2b",688 => x"c3a94590",689 => x"c45ae1d7",
690 => x"c50d1149",691 => x"c5bfd22f",692 => x"c67322ce",693 => x"c727016d",694 => x"c7db6c50",695 => x"c89061ba",696 => x"c945dfed",697 => x"c9fbe528",698 => x"cab26faa",699 => x"cb697db1",
700 => x"cc210d79",701 => x"ccd91d3e",702 => x"cd91ab39",703 => x"ce4ab5a3",704 => x"cf043ab3",705 => x"cfbe38a0",706 => x"d078ad9e",707 => x"d13397e2",708 => x"d1eef59f",709 => x"d2aac505",
710 => x"d3670446",711 => x"d423b191",712 => x"d4e0cb15",713 => x"d59e4eff",714 => x"d65c3b7c",715 => x"d71a8eb6",716 => x"d7d946d8",717 => x"d898620c",718 => x"d957de7b",719 => x"da17ba4b",
720 => x"dad7f3a3",721 => x"db9888a9",722 => x"dc597782",723 => x"dd1abe52",724 => x"dddc5b3b",725 => x"de9e4c61",726 => x"df608fe4",727 => x"e02323e6",728 => x"e0e60685",729 => x"e1a935e2",
730 => x"e26cb01b",731 => x"e330734d",732 => x"e3f47d96",733 => x"e4b8cd11",734 => x"e57d5fdb",735 => x"e642340e",736 => x"e70747c4",737 => x"e7cc9918",738 => x"e8922622",739 => x"e957ecfc",
740 => x"ea1debbc",741 => x"eae4207b",742 => x"ebaa894f",743 => x"ec712450",744 => x"ed37ef92",745 => x"edfee92c",746 => x"eec60f32",747 => x"ef8d5fb9",748 => x"f054d8d5",749 => x"f11c789b",
750 => x"f1e43d1d",751 => x"f2ac246e",752 => x"f3742ca2",753 => x"f43c53cb",754 => x"f50497fb",755 => x"f5ccf744",756 => x"f6956fb7",757 => x"f75dff66",758 => x"f826a462",759 => x"f8ef5cbc",
760 => x"f9b82684",761 => x"fa80ffcc",762 => x"fb49e6a3",763 => x"fc12d91a",764 => x"fcdbd542",765 => x"fda4d929",766 => x"fe6de2e1",767 => x"ff36f079",768 => x"00000000",769 => x"00c90f87",
770 => x"01921d1f",771 => x"025b26d7",772 => x"03242abe",773 => x"03ed26e6",774 => x"04b6195d",775 => x"057f0034",776 => x"0647d97c",777 => x"0710a344",778 => x"07d95b9e",779 => x"08a2009a",
780 => x"096a9049",781 => x"0a3308bc",782 => x"0afb6805",783 => x"0bc3ac35",784 => x"0c8bd35e",785 => x"0d53db92",786 => x"0e1bc2e3",787 => x"0ee38765",788 => x"0fab272b",789 => x"1072a047",
790 => x"1139f0ce",791 => x"120116d4",792 => x"12c8106e",793 => x"138edbb0",794 => x"145576b1",795 => x"151bdf85",796 => x"15e21444",797 => x"16a81304",798 => x"176dd9de",799 => x"183366e8",
800 => x"18f8b83c",801 => x"19bdcbf2",802 => x"1a82a025",803 => x"1b4732ef",804 => x"1c0b826a",805 => x"1ccf8cb3",806 => x"1d934fe5",807 => x"1e56ca1e",808 => x"1f19f97b",809 => x"1fdcdc1a",
810 => x"209f701c",811 => x"2161b39f",812 => x"2223a4c5",813 => x"22e541ae",814 => x"23a6887e",815 => x"24677757",816 => x"25280c5d",817 => x"25e845b5",818 => x"26a82185",819 => x"27679df4",
820 => x"2826b928",821 => x"28e5714a",822 => x"29a3c484",823 => x"2a61b101",824 => x"2b1f34eb",825 => x"2bdc4e6f",826 => x"2c98fbba",827 => x"2d553afb",828 => x"2e110a61",829 => x"2ecc681e",
830 => x"2f875262",831 => x"3041c760",832 => x"30fbc54d",833 => x"31b54a5d",834 => x"326e54c7",835 => x"3326e2c2",836 => x"33def287",837 => x"3496824f",838 => x"354d9056",839 => x"36041ad8",
840 => x"36ba2013",841 => x"376f9e46",842 => x"382493b0",843 => x"38d8fe93",844 => x"398cdd32",845 => x"3a402dd1",846 => x"3af2eeb7",847 => x"3ba51e29",848 => x"3c56ba70",849 => x"3d07c1d5",
850 => x"3db832a5",851 => x"3e680b2c",852 => x"3f1749b7",853 => x"3fc5ec97",854 => x"4073f21d",855 => x"4121589a",856 => x"41ce1e64",857 => x"427a41d0",858 => x"4325c135",859 => x"43d09aec",
860 => x"447acd50",861 => x"452456bc",862 => x"45cd358f",863 => x"46756827",864 => x"471cece6",865 => x"47c3c22e",866 => x"4869e664",867 => x"490f57ee",868 => x"49b41533",869 => x"4a581c9d",
870 => x"4afb6c97",871 => x"4b9e038f",872 => x"4c3fdff3",873 => x"4ce10034",874 => x"4d8162c4",875 => x"4e210617",876 => x"4ebfe8a4",877 => x"4f5e08e3",878 => x"4ffb654d",879 => x"5097fc5e",
880 => x"5133cc94",881 => x"51ced46e",882 => x"5269126e",883 => x"53028517",884 => x"539b2aef",885 => x"5433027d",886 => x"54ca0a4a",887 => x"556040e2",888 => x"55f5a4d2",889 => x"568a34a9",
890 => x"571deef9",891 => x"57b0d256",892 => x"5842dd54",893 => x"58d40e8c",894 => x"59646497",895 => x"59f3de12",896 => x"5a827999",897 => x"5b1035cf",898 => x"5b9d1153",899 => x"5c290acc",
900 => x"5cb420df",901 => x"5d3e5236",902 => x"5dc79d7c",903 => x"5e50015d",904 => x"5ed77c89",905 => x"5f5e0db3",906 => x"5fe3b38d",907 => x"60686cce",908 => x"60ec382f",909 => x"616f146b",
910 => x"61f1003e",911 => x"6271fa69",912 => x"62f201ac",913 => x"637114cc",914 => x"63ef328f",915 => x"646c59bf",916 => x"64e88926",917 => x"6563bf92",918 => x"65ddfbd3",919 => x"66573cbb",
920 => x"66cf811f",921 => x"6746c7d7",922 => x"67bd0fbc",923 => x"683257aa",924 => x"68a69e81",925 => x"6919e320",926 => x"698c246c",927 => x"69fd614a",928 => x"6a6d98a4",929 => x"6adcc964",
930 => x"6b4af278",931 => x"6bb812d0",932 => x"6c242960",933 => x"6c8f351c",934 => x"6cf934fb",935 => x"6d6227fa",936 => x"6dca0d14",937 => x"6e30e349",938 => x"6e96a99c",939 => x"6efb5f12",
940 => x"6f5f02b1",941 => x"6fc19385",942 => x"70231099",943 => x"708378fe",944 => x"70e2cbc6",945 => x"71410804",946 => x"719e2cd2",947 => x"71fa3948",948 => x"72552c84",949 => x"72af05a6",
950 => x"7307c3cf",951 => x"735f6626",952 => x"73b5ebd0",953 => x"740b53fa",954 => x"745f9dd0",955 => x"74b2c883",956 => x"7504d345",957 => x"7555bd4b",958 => x"75a585cf",959 => x"75f42c0a",
960 => x"7641af3c",961 => x"768e0ea5",962 => x"76d94988",963 => x"77235f2d",964 => x"776c4edb",965 => x"77b417df",966 => x"77fab988",967 => x"78403328",968 => x"78848413",969 => x"78c7aba1",
970 => x"7909a92c",971 => x"794a7c11",972 => x"798a23b1",973 => x"79c89f6d",974 => x"7a05eead",975 => x"7a4210d8",976 => x"7a7d055b",977 => x"7ab6cba3",978 => x"7aef6323",979 => x"7b26cb4f",
980 => x"7b5d039d",981 => x"7b920b89",982 => x"7bc5e28f",983 => x"7bf88830",984 => x"7c29fbee",985 => x"7c5a3d4f",986 => x"7c894bdd",987 => x"7cb72724",988 => x"7ce3ceb1",989 => x"7d0f4217",
990 => x"7d3980ec",991 => x"7d628ac5",992 => x"7d8a5f3f",993 => x"7db0fdf7",994 => x"7dd6668e",995 => x"7dfa98a7",996 => x"7e1d93e9",997 => x"7e3f57fe",998 => x"7e5fe493",999 => x"7e7f3956",
1000 => x"7e9d55fc",1001 => x"7eba3a39",1002 => x"7ed5e5c6",1003 => x"7ef0585f",1004 => x"7f0991c3",1005 => x"7f2191b3",1006 => x"7f3857f5",1007 => x"7f4de450",1008 => x"7f62368f",1009 => x"7f754e7f",
1010 => x"7f872bf2",1011 => x"7f97cebc",1012 => x"7fa736b4",1013 => x"7fb563b2",1014 => x"7fc25596",1015 => x"7fce0c3e",1016 => x"7fd8878d",1017 => x"7fe1c76b",1018 => x"7fe9cbbf",1019 => x"7ff09477",
1020 => x"7ff62182",1021 => x"7ffa72d1",1022 => x"7ffd8859",1023 => x"7fff6215");

constant TWIDDLE_FACTORS_IMAG : TWIDDLE_ARRAY(TWIDDLE_RANGE) := (0 => x"00000000",1 => x"ff36f079",2 => x"fe6de2e1",3 => x"fda4d929",4 => x"fcdbd542",5 => x"fc12d91a",6 => x"fb49e6a3",7 => x"fa80ffcc",8 => x"f9b82684",9 => x"f8ef5cbc",
10 => x"f826a462",11 => x"f75dff66",12 => x"f6956fb7",13 => x"f5ccf744",14 => x"f50497fb",15 => x"f43c53cb",16 => x"f3742ca2",17 => x"f2ac246e",18 => x"f1e43d1d",19 => x"f11c789b",
20 => x"f054d8d5",21 => x"ef8d5fb9",22 => x"eec60f32",23 => x"edfee92c",24 => x"ed37ef92",25 => x"ec712450",26 => x"ebaa894f",27 => x"eae4207b",28 => x"ea1debbc",29 => x"e957ecfc",
30 => x"e8922622",31 => x"e7cc9918",32 => x"e70747c4",33 => x"e642340e",34 => x"e57d5fdb",35 => x"e4b8cd11",36 => x"e3f47d96",37 => x"e330734d",38 => x"e26cb01b",39 => x"e1a935e2",
40 => x"e0e60685",41 => x"e02323e6",42 => x"df608fe4",43 => x"de9e4c61",44 => x"dddc5b3b",45 => x"dd1abe52",46 => x"dc597782",47 => x"db9888a9",48 => x"dad7f3a3",49 => x"da17ba4b",
50 => x"d957de7b",51 => x"d898620c",52 => x"d7d946d8",53 => x"d71a8eb6",54 => x"d65c3b7c",55 => x"d59e4eff",56 => x"d4e0cb15",57 => x"d423b191",58 => x"d3670446",59 => x"d2aac505",
60 => x"d1eef59f",61 => x"d13397e2",62 => x"d078ad9e",63 => x"cfbe38a0",64 => x"cf043ab3",65 => x"ce4ab5a3",66 => x"cd91ab39",67 => x"ccd91d3e",68 => x"cc210d79",69 => x"cb697db1",
70 => x"cab26faa",71 => x"c9fbe528",72 => x"c945dfed",73 => x"c89061ba",74 => x"c7db6c50",75 => x"c727016d",76 => x"c67322ce",77 => x"c5bfd22f",78 => x"c50d1149",79 => x"c45ae1d7",
80 => x"c3a94590",81 => x"c2f83e2b",82 => x"c247cd5b",83 => x"c197f4d4",84 => x"c0e8b649",85 => x"c03a1369",86 => x"bf8c0de3",87 => x"bedea766",88 => x"be31e19c",89 => x"bd85be30",
90 => x"bcda3ecb",91 => x"bc2f6514",92 => x"bb8532b0",93 => x"badba944",94 => x"ba32ca71",95 => x"b98a97d9",96 => x"b8e3131a",97 => x"b83c3dd2",98 => x"b796199c",99 => x"b6f0a812",
100 => x"b64beacd",101 => x"b5a7e363",102 => x"b5049369",103 => x"b461fc71",104 => x"b3c0200d",105 => x"b31effcc",106 => x"b27e9d3c",107 => x"b1def9e9",108 => x"b140175c",109 => x"b0a1f71d",
110 => x"b0049ab3",111 => x"af6803a2",112 => x"aecc336c",113 => x"ae312b92",114 => x"ad96ed92",115 => x"acfd7ae9",116 => x"ac64d511",117 => x"abccfd83",118 => x"ab35f5b6",119 => x"aa9fbf1e",
120 => x"aa0a5b2e",121 => x"a975cb57",122 => x"a8e21107",123 => x"a84f2daa",124 => x"a7bd22ac",125 => x"a72bf174",126 => x"a69b9b69",127 => x"a60c21ee",128 => x"a57d8667",129 => x"a4efca31",
130 => x"a462eead",131 => x"a3d6f534",132 => x"a34bdf21",133 => x"a2c1adca",134 => x"a2386284",135 => x"a1affea3",136 => x"a1288377",137 => x"a0a1f24d",138 => x"a01c4c73",139 => x"9f979332",
140 => x"9f13c7d1",141 => x"9e90eb95",142 => x"9e0effc2",143 => x"9d8e0597",144 => x"9d0dfe54",145 => x"9c8eeb34",146 => x"9c10cd71",147 => x"9b93a641",148 => x"9b1776da",149 => x"9a9c406e",
150 => x"9a22042d",151 => x"99a8c345",152 => x"99307ee1",153 => x"98b93829",154 => x"9842f044",155 => x"97cda856",156 => x"9759617f",157 => x"96e61ce0",158 => x"9673db94",159 => x"96029eb6",
160 => x"9592675c",161 => x"9523369c",162 => x"94b50d88",163 => x"9447ed30",164 => x"93dbd6a0",165 => x"9370cae4",166 => x"9306cb05",167 => x"929dd806",168 => x"9235f2ec",169 => x"91cf1cb7",
170 => x"91695664",171 => x"9104a0ee",172 => x"90a0fd4f",173 => x"903e6c7b",174 => x"8fdcef67",175 => x"8f7c8702",176 => x"8f1d343a",177 => x"8ebef7fc",178 => x"8e61d32e",179 => x"8e05c6b8",
180 => x"8daad37c",181 => x"8d50fa5a",182 => x"8cf83c31",183 => x"8ca099da",184 => x"8c4a1430",185 => x"8bf4ac06",186 => x"8ba06230",187 => x"8b4d377d",188 => x"8afb2cbb",189 => x"8aaa42b5",
190 => x"8a5a7a31",191 => x"8a0bd3f6",192 => x"89be50c4",193 => x"8971f15b",194 => x"8926b678",195 => x"88dca0d3",196 => x"8893b125",197 => x"884be821",198 => x"88054678",199 => x"87bfccd8",
200 => x"877b7bed",201 => x"8738545f",202 => x"86f656d4",203 => x"86b583ef",204 => x"8675dc4f",205 => x"86376093",206 => x"85fa1153",207 => x"85bdef28",208 => x"8582faa5",209 => x"8549345d",
210 => x"85109cdd",211 => x"84d934b1",212 => x"84a2fc63",213 => x"846df477",214 => x"843a1d71",215 => x"840777d0",216 => x"83d60412",217 => x"83a5c2b1",218 => x"8376b423",219 => x"8348d8dc",
220 => x"831c314f",221 => x"82f0bde9",222 => x"82c67f14",223 => x"829d753b",224 => x"8275a0c1",225 => x"824f0209",226 => x"82299972",227 => x"82056759",228 => x"81e26c17",229 => x"81c0a802",
230 => x"81a01b6d",231 => x"8180c6aa",232 => x"8162aa04",233 => x"8145c5c7",234 => x"812a1a3a",235 => x"810fa7a1",236 => x"80f66e3d",237 => x"80de6e4d",238 => x"80c7a80b",239 => x"80b21bb0",
240 => x"809dc971",241 => x"808ab181",242 => x"8078d40e",243 => x"80683144",244 => x"8058c94c",245 => x"804a9c4e",246 => x"803daa6a",247 => x"8031f3c2",248 => x"80277873",249 => x"801e3895",
250 => x"80163441",251 => x"800f6b89",252 => x"8009de7e",253 => x"80058d2f",254 => x"800277a6",255 => x"80009dea",256 => x"80000000",257 => x"80009dea",258 => x"800277a6",259 => x"80058d2f",
260 => x"8009de7e",261 => x"800f6b89",262 => x"80163441",263 => x"801e3895",264 => x"80277873",265 => x"8031f3c2",266 => x"803daa6a",267 => x"804a9c4e",268 => x"8058c94c",269 => x"80683144",
270 => x"8078d40e",271 => x"808ab181",272 => x"809dc971",273 => x"80b21bb0",274 => x"80c7a80b",275 => x"80de6e4d",276 => x"80f66e3d",277 => x"810fa7a1",278 => x"812a1a3a",279 => x"8145c5c7",
280 => x"8162aa04",281 => x"8180c6aa",282 => x"81a01b6d",283 => x"81c0a802",284 => x"81e26c17",285 => x"82056759",286 => x"82299972",287 => x"824f0209",288 => x"8275a0c1",289 => x"829d753b",
290 => x"82c67f14",291 => x"82f0bde9",292 => x"831c314f",293 => x"8348d8dc",294 => x"8376b423",295 => x"83a5c2b1",296 => x"83d60412",297 => x"840777d0",298 => x"843a1d71",299 => x"846df477",
300 => x"84a2fc63",301 => x"84d934b1",302 => x"85109cdd",303 => x"8549345d",304 => x"8582faa5",305 => x"85bdef28",306 => x"85fa1153",307 => x"86376093",308 => x"8675dc4f",309 => x"86b583ef",
310 => x"86f656d4",311 => x"8738545f",312 => x"877b7bed",313 => x"87bfccd8",314 => x"88054678",315 => x"884be821",316 => x"8893b125",317 => x"88dca0d3",318 => x"8926b678",319 => x"8971f15b",
320 => x"89be50c4",321 => x"8a0bd3f6",322 => x"8a5a7a31",323 => x"8aaa42b5",324 => x"8afb2cbb",325 => x"8b4d377d",326 => x"8ba06230",327 => x"8bf4ac06",328 => x"8c4a1430",329 => x"8ca099da",
330 => x"8cf83c31",331 => x"8d50fa5a",332 => x"8daad37c",333 => x"8e05c6b8",334 => x"8e61d32e",335 => x"8ebef7fc",336 => x"8f1d343a",337 => x"8f7c8702",338 => x"8fdcef67",339 => x"903e6c7b",
340 => x"90a0fd4f",341 => x"9104a0ee",342 => x"91695664",343 => x"91cf1cb7",344 => x"9235f2ec",345 => x"929dd806",346 => x"9306cb05",347 => x"9370cae4",348 => x"93dbd6a0",349 => x"9447ed30",
350 => x"94b50d88",351 => x"9523369c",352 => x"9592675c",353 => x"96029eb6",354 => x"9673db94",355 => x"96e61ce0",356 => x"9759617f",357 => x"97cda856",358 => x"9842f044",359 => x"98b93829",
360 => x"99307ee1",361 => x"99a8c345",362 => x"9a22042d",363 => x"9a9c406e",364 => x"9b1776da",365 => x"9b93a641",366 => x"9c10cd71",367 => x"9c8eeb34",368 => x"9d0dfe54",369 => x"9d8e0597",
370 => x"9e0effc2",371 => x"9e90eb95",372 => x"9f13c7d1",373 => x"9f979332",374 => x"a01c4c73",375 => x"a0a1f24d",376 => x"a1288377",377 => x"a1affea3",378 => x"a2386284",379 => x"a2c1adca",
380 => x"a34bdf21",381 => x"a3d6f534",382 => x"a462eead",383 => x"a4efca31",384 => x"a57d8667",385 => x"a60c21ee",386 => x"a69b9b69",387 => x"a72bf174",388 => x"a7bd22ac",389 => x"a84f2daa",
390 => x"a8e21107",391 => x"a975cb57",392 => x"aa0a5b2e",393 => x"aa9fbf1e",394 => x"ab35f5b6",395 => x"abccfd83",396 => x"ac64d511",397 => x"acfd7ae9",398 => x"ad96ed92",399 => x"ae312b92",
400 => x"aecc336c",401 => x"af6803a2",402 => x"b0049ab3",403 => x"b0a1f71d",404 => x"b140175c",405 => x"b1def9e9",406 => x"b27e9d3c",407 => x"b31effcc",408 => x"b3c0200d",409 => x"b461fc71",
410 => x"b5049369",411 => x"b5a7e363",412 => x"b64beacd",413 => x"b6f0a812",414 => x"b796199c",415 => x"b83c3dd2",416 => x"b8e3131a",417 => x"b98a97d9",418 => x"ba32ca71",419 => x"badba944",
420 => x"bb8532b0",421 => x"bc2f6514",422 => x"bcda3ecb",423 => x"bd85be30",424 => x"be31e19c",425 => x"bedea766",426 => x"bf8c0de3",427 => x"c03a1369",428 => x"c0e8b649",429 => x"c197f4d4",
430 => x"c247cd5b",431 => x"c2f83e2b",432 => x"c3a94590",433 => x"c45ae1d7",434 => x"c50d1149",435 => x"c5bfd22f",436 => x"c67322ce",437 => x"c727016d",438 => x"c7db6c50",439 => x"c89061ba",
440 => x"c945dfed",441 => x"c9fbe528",442 => x"cab26faa",443 => x"cb697db1",444 => x"cc210d79",445 => x"ccd91d3e",446 => x"cd91ab39",447 => x"ce4ab5a3",448 => x"cf043ab3",449 => x"cfbe38a0",
450 => x"d078ad9e",451 => x"d13397e2",452 => x"d1eef59f",453 => x"d2aac505",454 => x"d3670446",455 => x"d423b191",456 => x"d4e0cb15",457 => x"d59e4eff",458 => x"d65c3b7c",459 => x"d71a8eb6",
460 => x"d7d946d8",461 => x"d898620c",462 => x"d957de7b",463 => x"da17ba4b",464 => x"dad7f3a3",465 => x"db9888a9",466 => x"dc597782",467 => x"dd1abe52",468 => x"dddc5b3b",469 => x"de9e4c61",
470 => x"df608fe4",471 => x"e02323e6",472 => x"e0e60685",473 => x"e1a935e2",474 => x"e26cb01b",475 => x"e330734d",476 => x"e3f47d96",477 => x"e4b8cd11",478 => x"e57d5fdb",479 => x"e642340e",
480 => x"e70747c4",481 => x"e7cc9918",482 => x"e8922622",483 => x"e957ecfc",484 => x"ea1debbc",485 => x"eae4207b",486 => x"ebaa894f",487 => x"ec712450",488 => x"ed37ef92",489 => x"edfee92c",
490 => x"eec60f32",491 => x"ef8d5fb9",492 => x"f054d8d5",493 => x"f11c789b",494 => x"f1e43d1d",495 => x"f2ac246e",496 => x"f3742ca2",497 => x"f43c53cb",498 => x"f50497fb",499 => x"f5ccf744",
500 => x"f6956fb7",501 => x"f75dff66",502 => x"f826a462",503 => x"f8ef5cbc",504 => x"f9b82684",505 => x"fa80ffcc",506 => x"fb49e6a3",507 => x"fc12d91a",508 => x"fcdbd542",509 => x"fda4d929",
510 => x"fe6de2e1",511 => x"ff36f079",512 => x"00000000",513 => x"00c90f87",514 => x"01921d1f",515 => x"025b26d7",516 => x"03242abe",517 => x"03ed26e6",518 => x"04b6195d",519 => x"057f0034",
520 => x"0647d97c",521 => x"0710a344",522 => x"07d95b9e",523 => x"08a2009a",524 => x"096a9049",525 => x"0a3308bc",526 => x"0afb6805",527 => x"0bc3ac35",528 => x"0c8bd35e",529 => x"0d53db92",
530 => x"0e1bc2e3",531 => x"0ee38765",532 => x"0fab272b",533 => x"1072a047",534 => x"1139f0ce",535 => x"120116d4",536 => x"12c8106e",537 => x"138edbb0",538 => x"145576b1",539 => x"151bdf85",
540 => x"15e21444",541 => x"16a81304",542 => x"176dd9de",543 => x"183366e8",544 => x"18f8b83c",545 => x"19bdcbf2",546 => x"1a82a025",547 => x"1b4732ef",548 => x"1c0b826a",549 => x"1ccf8cb3",
550 => x"1d934fe5",551 => x"1e56ca1e",552 => x"1f19f97b",553 => x"1fdcdc1a",554 => x"209f701c",555 => x"2161b39f",556 => x"2223a4c5",557 => x"22e541ae",558 => x"23a6887e",559 => x"24677757",
560 => x"25280c5d",561 => x"25e845b5",562 => x"26a82185",563 => x"27679df4",564 => x"2826b928",565 => x"28e5714a",566 => x"29a3c484",567 => x"2a61b101",568 => x"2b1f34eb",569 => x"2bdc4e6f",
570 => x"2c98fbba",571 => x"2d553afb",572 => x"2e110a61",573 => x"2ecc681e",574 => x"2f875262",575 => x"3041c760",576 => x"30fbc54d",577 => x"31b54a5d",578 => x"326e54c7",579 => x"3326e2c2",
580 => x"33def287",581 => x"3496824f",582 => x"354d9056",583 => x"36041ad8",584 => x"36ba2013",585 => x"376f9e46",586 => x"382493b0",587 => x"38d8fe93",588 => x"398cdd32",589 => x"3a402dd1",
590 => x"3af2eeb7",591 => x"3ba51e29",592 => x"3c56ba70",593 => x"3d07c1d5",594 => x"3db832a5",595 => x"3e680b2c",596 => x"3f1749b7",597 => x"3fc5ec97",598 => x"4073f21d",599 => x"4121589a",
600 => x"41ce1e64",601 => x"427a41d0",602 => x"4325c135",603 => x"43d09aec",604 => x"447acd50",605 => x"452456bc",606 => x"45cd358f",607 => x"46756827",608 => x"471cece6",609 => x"47c3c22e",
610 => x"4869e664",611 => x"490f57ee",612 => x"49b41533",613 => x"4a581c9d",614 => x"4afb6c97",615 => x"4b9e038f",616 => x"4c3fdff3",617 => x"4ce10034",618 => x"4d8162c4",619 => x"4e210617",
620 => x"4ebfe8a4",621 => x"4f5e08e3",622 => x"4ffb654d",623 => x"5097fc5e",624 => x"5133cc94",625 => x"51ced46e",626 => x"5269126e",627 => x"53028517",628 => x"539b2aef",629 => x"5433027d",
630 => x"54ca0a4a",631 => x"556040e2",632 => x"55f5a4d2",633 => x"568a34a9",634 => x"571deef9",635 => x"57b0d256",636 => x"5842dd54",637 => x"58d40e8c",638 => x"59646497",639 => x"59f3de12",
640 => x"5a827999",641 => x"5b1035cf",642 => x"5b9d1153",643 => x"5c290acc",644 => x"5cb420df",645 => x"5d3e5236",646 => x"5dc79d7c",647 => x"5e50015d",648 => x"5ed77c89",649 => x"5f5e0db3",
650 => x"5fe3b38d",651 => x"60686cce",652 => x"60ec382f",653 => x"616f146b",654 => x"61f1003e",655 => x"6271fa69",656 => x"62f201ac",657 => x"637114cc",658 => x"63ef328f",659 => x"646c59bf",
660 => x"64e88926",661 => x"6563bf92",662 => x"65ddfbd3",663 => x"66573cbb",664 => x"66cf811f",665 => x"6746c7d7",666 => x"67bd0fbc",667 => x"683257aa",668 => x"68a69e81",669 => x"6919e320",
670 => x"698c246c",671 => x"69fd614a",672 => x"6a6d98a4",673 => x"6adcc964",674 => x"6b4af278",675 => x"6bb812d0",676 => x"6c242960",677 => x"6c8f351c",678 => x"6cf934fb",679 => x"6d6227fa",
680 => x"6dca0d14",681 => x"6e30e349",682 => x"6e96a99c",683 => x"6efb5f12",684 => x"6f5f02b1",685 => x"6fc19385",686 => x"70231099",687 => x"708378fe",688 => x"70e2cbc6",689 => x"71410804",
690 => x"719e2cd2",691 => x"71fa3948",692 => x"72552c84",693 => x"72af05a6",694 => x"7307c3cf",695 => x"735f6626",696 => x"73b5ebd0",697 => x"740b53fa",698 => x"745f9dd0",699 => x"74b2c883",
700 => x"7504d345",701 => x"7555bd4b",702 => x"75a585cf",703 => x"75f42c0a",704 => x"7641af3c",705 => x"768e0ea5",706 => x"76d94988",707 => x"77235f2d",708 => x"776c4edb",709 => x"77b417df",
710 => x"77fab988",711 => x"78403328",712 => x"78848413",713 => x"78c7aba1",714 => x"7909a92c",715 => x"794a7c11",716 => x"798a23b1",717 => x"79c89f6d",718 => x"7a05eead",719 => x"7a4210d8",
720 => x"7a7d055b",721 => x"7ab6cba3",722 => x"7aef6323",723 => x"7b26cb4f",724 => x"7b5d039d",725 => x"7b920b89",726 => x"7bc5e28f",727 => x"7bf88830",728 => x"7c29fbee",729 => x"7c5a3d4f",
730 => x"7c894bdd",731 => x"7cb72724",732 => x"7ce3ceb1",733 => x"7d0f4217",734 => x"7d3980ec",735 => x"7d628ac5",736 => x"7d8a5f3f",737 => x"7db0fdf7",738 => x"7dd6668e",739 => x"7dfa98a7",
740 => x"7e1d93e9",741 => x"7e3f57fe",742 => x"7e5fe493",743 => x"7e7f3956",744 => x"7e9d55fc",745 => x"7eba3a39",746 => x"7ed5e5c6",747 => x"7ef0585f",748 => x"7f0991c3",749 => x"7f2191b3",
750 => x"7f3857f5",751 => x"7f4de450",752 => x"7f62368f",753 => x"7f754e7f",754 => x"7f872bf2",755 => x"7f97cebc",756 => x"7fa736b4",757 => x"7fb563b2",758 => x"7fc25596",759 => x"7fce0c3e",
760 => x"7fd8878d",761 => x"7fe1c76b",762 => x"7fe9cbbf",763 => x"7ff09477",764 => x"7ff62182",765 => x"7ffa72d1",766 => x"7ffd8859",767 => x"7fff6215",768 => x"7fffffff",769 => x"7fff6215",
770 => x"7ffd8859",771 => x"7ffa72d1",772 => x"7ff62182",773 => x"7ff09477",774 => x"7fe9cbbf",775 => x"7fe1c76b",776 => x"7fd8878d",777 => x"7fce0c3e",778 => x"7fc25596",779 => x"7fb563b2",
780 => x"7fa736b4",781 => x"7f97cebc",782 => x"7f872bf2",783 => x"7f754e7f",784 => x"7f62368f",785 => x"7f4de450",786 => x"7f3857f5",787 => x"7f2191b3",788 => x"7f0991c3",789 => x"7ef0585f",
790 => x"7ed5e5c6",791 => x"7eba3a39",792 => x"7e9d55fc",793 => x"7e7f3956",794 => x"7e5fe493",795 => x"7e3f57fe",796 => x"7e1d93e9",797 => x"7dfa98a7",798 => x"7dd6668e",799 => x"7db0fdf7",
800 => x"7d8a5f3f",801 => x"7d628ac5",802 => x"7d3980ec",803 => x"7d0f4217",804 => x"7ce3ceb1",805 => x"7cb72724",806 => x"7c894bdd",807 => x"7c5a3d4f",808 => x"7c29fbee",809 => x"7bf88830",
810 => x"7bc5e28f",811 => x"7b920b89",812 => x"7b5d039d",813 => x"7b26cb4f",814 => x"7aef6323",815 => x"7ab6cba3",816 => x"7a7d055b",817 => x"7a4210d8",818 => x"7a05eead",819 => x"79c89f6d",
820 => x"798a23b1",821 => x"794a7c11",822 => x"7909a92c",823 => x"78c7aba1",824 => x"78848413",825 => x"78403328",826 => x"77fab988",827 => x"77b417df",828 => x"776c4edb",829 => x"77235f2d",
830 => x"76d94988",831 => x"768e0ea5",832 => x"7641af3c",833 => x"75f42c0a",834 => x"75a585cf",835 => x"7555bd4b",836 => x"7504d345",837 => x"74b2c883",838 => x"745f9dd0",839 => x"740b53fa",
840 => x"73b5ebd0",841 => x"735f6626",842 => x"7307c3cf",843 => x"72af05a6",844 => x"72552c84",845 => x"71fa3948",846 => x"719e2cd2",847 => x"71410804",848 => x"70e2cbc6",849 => x"708378fe",
850 => x"70231099",851 => x"6fc19385",852 => x"6f5f02b1",853 => x"6efb5f12",854 => x"6e96a99c",855 => x"6e30e349",856 => x"6dca0d14",857 => x"6d6227fa",858 => x"6cf934fb",859 => x"6c8f351c",
860 => x"6c242960",861 => x"6bb812d0",862 => x"6b4af278",863 => x"6adcc964",864 => x"6a6d98a4",865 => x"69fd614a",866 => x"698c246c",867 => x"6919e320",868 => x"68a69e81",869 => x"683257aa",
870 => x"67bd0fbc",871 => x"6746c7d7",872 => x"66cf811f",873 => x"66573cbb",874 => x"65ddfbd3",875 => x"6563bf92",876 => x"64e88926",877 => x"646c59bf",878 => x"63ef328f",879 => x"637114cc",
880 => x"62f201ac",881 => x"6271fa69",882 => x"61f1003e",883 => x"616f146b",884 => x"60ec382f",885 => x"60686cce",886 => x"5fe3b38d",887 => x"5f5e0db3",888 => x"5ed77c89",889 => x"5e50015d",
890 => x"5dc79d7c",891 => x"5d3e5236",892 => x"5cb420df",893 => x"5c290acc",894 => x"5b9d1153",895 => x"5b1035cf",896 => x"5a827999",897 => x"59f3de12",898 => x"59646497",899 => x"58d40e8c",
900 => x"5842dd54",901 => x"57b0d256",902 => x"571deef9",903 => x"568a34a9",904 => x"55f5a4d2",905 => x"556040e2",906 => x"54ca0a4a",907 => x"5433027d",908 => x"539b2aef",909 => x"53028517",
910 => x"5269126e",911 => x"51ced46e",912 => x"5133cc94",913 => x"5097fc5e",914 => x"4ffb654d",915 => x"4f5e08e3",916 => x"4ebfe8a4",917 => x"4e210617",918 => x"4d8162c4",919 => x"4ce10034",
920 => x"4c3fdff3",921 => x"4b9e038f",922 => x"4afb6c97",923 => x"4a581c9d",924 => x"49b41533",925 => x"490f57ee",926 => x"4869e664",927 => x"47c3c22e",928 => x"471cece6",929 => x"46756827",
930 => x"45cd358f",931 => x"452456bc",932 => x"447acd50",933 => x"43d09aec",934 => x"4325c135",935 => x"427a41d0",936 => x"41ce1e64",937 => x"4121589a",938 => x"4073f21d",939 => x"3fc5ec97",
940 => x"3f1749b7",941 => x"3e680b2c",942 => x"3db832a5",943 => x"3d07c1d5",944 => x"3c56ba70",945 => x"3ba51e29",946 => x"3af2eeb7",947 => x"3a402dd1",948 => x"398cdd32",949 => x"38d8fe93",
950 => x"382493b0",951 => x"376f9e46",952 => x"36ba2013",953 => x"36041ad8",954 => x"354d9056",955 => x"3496824f",956 => x"33def287",957 => x"3326e2c2",958 => x"326e54c7",959 => x"31b54a5d",
960 => x"30fbc54d",961 => x"3041c760",962 => x"2f875262",963 => x"2ecc681e",964 => x"2e110a61",965 => x"2d553afb",966 => x"2c98fbba",967 => x"2bdc4e6f",968 => x"2b1f34eb",969 => x"2a61b101",
970 => x"29a3c484",971 => x"28e5714a",972 => x"2826b928",973 => x"27679df4",974 => x"26a82185",975 => x"25e845b5",976 => x"25280c5d",977 => x"24677757",978 => x"23a6887e",979 => x"22e541ae",
980 => x"2223a4c5",981 => x"2161b39f",982 => x"209f701c",983 => x"1fdcdc1a",984 => x"1f19f97b",985 => x"1e56ca1e",986 => x"1d934fe5",987 => x"1ccf8cb3",988 => x"1c0b826a",989 => x"1b4732ef",
990 => x"1a82a025",991 => x"19bdcbf2",992 => x"18f8b83c",993 => x"183366e8",994 => x"176dd9de",995 => x"16a81304",996 => x"15e21444",997 => x"151bdf85",998 => x"145576b1",999 => x"138edbb0",
1000 => x"12c8106e",1001 => x"120116d4",1002 => x"1139f0ce",1003 => x"1072a047",1004 => x"0fab272b",1005 => x"0ee38765",1006 => x"0e1bc2e3",1007 => x"0d53db92",1008 => x"0c8bd35e",1009 => x"0bc3ac35",
1010 => x"0afb6805",1011 => x"0a3308bc",1012 => x"096a9049",1013 => x"08a2009a",1014 => x"07d95b9e",1015 => x"0710a344",1016 => x"0647d97c",1017 => x"057f0034",1018 => x"04b6195d",1019 => x"03ed26e6",
1020 => x"03242abe",1021 => x"025b26d7",1022 => x"01921d1f",1023 => x"00c90f87");

constant ZERO : std_logic_vector(DATA_RANGE) := (others => '0');

constant NEGATIVE_ONE : std_logic_vector(DATA_RANGE) := ((DATA_WIDTH - 1) => '1', others => '0');

end user_pkg;